//module procesador(
//	input clk;
//	input rst;
//	input test;
//	
//	input btn_back,
//	input btn_next,
//	input btn_comer_inc,     		   
//	input btn_curar_dec,				
//	input sns_prox,
//	input sns_temp,
//	input sns_luz,

//	input inSalud,
//	input inAnimo,
//	input inComida,
//	input inEnergia,
//	input inState,
//	input inDias,
//);
//
////	reg [2:0] SALUD;     			 
////	reg [2:0] ANIMO;      
////	reg [2:0] COMIDA;     
////	reg [2:0] ENERGIA;
////	reg [3:0] STATE;					
////	reg [5:0] DIAS;      			
////	reg [2:0] reg_stat;   			
////	reg [31:0] second_counter;		
////	reg [31:0] minute_counter;  	
////	reg time_enable;
//
////	initial begin
////		SALUD   = 3'd5;
////		ANIMO   = 3'd5;
////		COMIDA  = 3'd5;
////		ENERGIA = 3'd5;
////		DIAS    = 6'd0;
////		STATE   = 4'b1111;
////		reg_stat = 3'd0;
////		second_counter = 32'd0;
////		minute_counter = 32'd0;
////		time_enable <= 1'b0;
////	end
//
//	wire wire_clk_div;
//
//	divisor div1(
//		.clkd(clk),
//		.clk2(wire_clk_div)
//	);
//
//	always @(posedge (wire_clk_div)) begin
//	
//		if (rst == 0) begin
//
////			SALUD   	 <= 3'd5;
////			ANIMO   	 <= 3'd5;
////			COMIDA  	 <= 3'd5;
////			ENERGIA 	 <= 3'd5;
////			DIAS	 	 <= 6'd0;
////			STATE		 <= 4'd15;
////			second_counter = 32'd0;
////			minute_counter = 32'd0;
////			time_enable <= 1'd0;
//
//		end else begin
//		
//		if (SALUD < 3'd2 && STATE[3] == 1'b1) begin
//			STATE <= {1'b0, STATE[2:0]}; 
//		end else if (SALUD >= 3'd2 && STATE[3] == 1'b0) begin
//			STATE <= {1'b1, STATE[2:0]};
//		end
//		
//		if (ANIMO < 3'd2 && STATE[2] == 1'b1) begin
//			STATE <= {STATE[3], 1'b0, STATE[1:0]}; 
//		end else if (ANIMO >= 3'd2 && STATE[2] == 1'b0) begin
//			STATE <= {STATE[3], 1'b1, STATE[1:0]};
//		end
//		
//		if (COMIDA < 3'd2 && STATE[1] == 1'b1) begin
//			STATE <= {STATE[3:2], 1'b0, STATE[0]}; 
//		end else if (COMIDA >= 3'd2 && STATE[1] == 1'b0) begin
//			STATE <= {STATE[3:2], 1'b1, STATE[0]};
//		end
//		
//		if (ENERGIA < 3'd2 && STATE[0] == 1'b1) begin
//			STATE <= {STATE[3:1],1'b0}; 
//		end else if (ENERGIA >= 3'd2 && STATE[0] == 1'b0) begin
//			STATE <= {STATE[3:1], 1'b1};
//		end
//
//		if (time_enable) begin
//				
//				if (second_counter < wire_clk_div * (10)) begin // 5*(tiempo_cambio) = multiplicador; 5 => 60s_divisor/12s_reales
//					
//					second_counter <= second_counter + 1;
//				
//				end else begin
//				
//					second_counter <= 32'd0;      // Reiniciar el contador de segundos
//					minute_counter <= minute_counter + 1;  // Incrementar los minutos
//
//					if (second_counter >= MINUTES_TO_INCREMENT_DAYS) begin
////					if (minute_counter >= MINUTES_TO_INCREMENT_DAYS) begin
//						minute_counter <= 32'd0;  
//						DIAS <= DIAS + 1;         
//
//						if (DIAS >= 6'd32) begin
//
//							SALUD			<= 3'd0;
//							ANIMO			<= 3'd0;
//							COMIDA		<= 3'd0;
//							ENERGIA		<= 3'd0;
//							DIAS			<= 6'd0;
//							STATE			<= 4'd0;
//							time_enable <= 1'd0;
//						
//						end
//					end
//				end
//			end
//
//			if (btn_next == 0) begin
//				reg_stat <= (reg_stat < 3'd5) ? reg_stat + 1 : 3'd0;
//			end
//
//			if (btn_back == 0) begin
//				reg_stat <= (reg_stat > 3'd0) ? reg_stat - 1 : 3'd5;
//			end
//			
//			if (btn_comer_inc == 0) begin
//				
//				case (reg_stat)														
//					
//					3'd0: SALUD   <= (SALUD < 3'd5)   ? SALUD + 1   : SALUD;			
//					3'd1: ANIMO   <= (ANIMO < 3'd5)   ? ANIMO + 1   : ANIMO;			
//					3'd2: COMIDA  <= (COMIDA < 3'd5)  ? COMIDA + 1  : COMIDA;		
//					3'd3: ENERGIA <= (ENERGIA < 3'd5) ? ENERGIA + 1 : ENERGIA;	
//					3'd4: begin
//								DIAS    <= (DIAS < 6'd32)   ? DIAS + 1 : 6'd0;
//								SALUD   <= (DIAS >= 6'd32)  ? 4'd0     : SALUD;
//								ANIMO   <= (DIAS >= 6'd32)  ? 4'd0     : ANIMO;
//								COMIDA  <= (DIAS >= 6'd32)  ? 4'd0     : COMIDA;
//								ENERGIA <= (DIAS >= 6'd32)  ? 4'd0     : ENERGIA;
//								STATE   <= (DIAS >= 6'd32)  ? 4'd0     : STATE;
//							end
//					3'd5: STATE   <= (STATE < 4'd15)  ? STATE + 1   : STATE;
//
//				endcase
//				
//			end
//
//			if (btn_curar_dec == 0) begin
//				
//				case (reg_stat)	
//				
//					3'd0: if (SALUD > 3'd0) SALUD <= SALUD - 1;			
//					3'd1: if (ANIMO > 3'd0) ANIMO <= ANIMO - 1;			
//					3'd2: if (COMIDA > 3'd0) COMIDA <= COMIDA - 1;		
//					3'd3: if (ENERGIA > 3'd0) ENERGIA <= ENERGIA - 1;	
//					3'd4: if (DIAS > 6'd0) DIAS <= DIAS - 1;
//					3'd5: if (STATE > 4'd0) STATE <= STATE - 1;	
//									
//				endcase
//				
//			end
//
//			case (reg_stat)
//
//				3'd0: begin
//					stat_name <= 4'd5;     
//					stat_value <= SALUD;
//					state <= STATE;
//				end
//
//				3'd1: begin
//					stat_name <= 4'ha;     
//					stat_value <= ANIMO;
//					state <= STATE;   
//				end
//
//				3'd2: begin
//					stat_name <= 4'hc;     
//					stat_value <= COMIDA;
//					state <= STATE;  
//				end
//
//				3'd3: begin
//					stat_name <= 4'he;     
//					stat_value <= ENERGIA;
//					state <= STATE; 
//				end
//
//				3'd4: begin
//					stat_name <= 4'hd;     
//					stat_value <= DIAS[5:0];
//					state <= STATE; 
//				end
//				
//				3'd5: begin
//					stat_name <= 4'hf;     
//					stat_value <= STATE;   
//				end
//
//			endcase
//			
//		end
//		
//	end
//	
//endmodule