module spi_master #(parameter DATA_SIZE = 9)(
    input wire clk,
    input wire rst,
    input wire [DATA_SIZE-1:0] input_data,
    input wire available_data,
    output wire spi_sck,
    output reg spi_mosi,
    output reg spi_dc,
    output wire spi_cs,
    output reg idle
);

reg [0:2] data_bit_counter = 3'b0;
reg [DATA_SIZE-1:0] data_reg;
reg sck_reg;
reg cs_reg;

initial begin
    sck_reg <= 1'b1;
    data_reg <= 1'b0;
    data_bit_counter <= 3'b0;
    idle <= 1'b1;
    cs_reg <= 1'b0;
    spi_mosi <= 1'b0;
    spi_dc <= 1'b1;
end

wire dc = data_reg[8];
wire [0:DATA_SIZE-2] real_data = data_reg[DATA_SIZE-2:0];

assign spi_sck = sck_reg & cs_reg;
assign spi_cs = !cs_reg;

always @(posedge clk or posedge rst) begin
    if (rst) begin
        sck_reg <= 1'b1;
        data_reg <= 1'b0;
        data_bit_counter <= 3'b0;
        idle <= 1'b1;
        cs_reg <= 1'b0;
        spi_mosi <= 1'b0;
        spi_dc <= 1'b1;
    end else begin
        if (available_data) begin
            data_reg <= input_data;
            idle <= 1'b0;
            data_bit_counter <= 3'b0;
            cs_reg <= 1'b1; // Assert CS when starting data transfer
        end
        if (!idle) begin
            sck_reg <= !sck_reg;
            if (sck_reg) begin
                spi_dc <= dc;
                spi_mosi <= real_data[data_bit_counter];
                data_bit_counter <= data_bit_counter + 1'b1;
                if (data_bit_counter == (DATA_SIZE-1)) begin
                    idle <= 1'b1; // Set idle after completing data transfer
                end
            end
        end else begin
            sck_reg <= 1'b1;
            if (sck_reg) begin
                cs_reg <= 1'b0; // Deassert CS when idle
                spi_dc <= 1'b1;
            end
        end
    end
end
endmodule